module hello;
	initial begin
		$display("hello.");
		$finish;
	end
endmodule
